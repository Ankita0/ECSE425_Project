LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_signed.all;

ENTITY IF_mux_behaviour IS

PORT(
IN;
IN;
OUT);
END IF_mux_behaviour;


ARCHITECTURE mux_behaviour IS


END mux_behaviour;