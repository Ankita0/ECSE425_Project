library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity execute_stage is


end execute_stage;


architecture testbed of execute_stage is

begin



end testbed;
