library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity execute_stage is

	Port(A,B,C,D,E: in std_logic_vector (31 downto 0)
			W,X,Y.Z: out std_logic_vector(31 downto 0));


end execute_stage;


architecture testbed of execute_stage is

begin



end testbed;
