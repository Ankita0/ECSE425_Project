library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY Zero is 

PORT();

end Zero;


Architecture arch of zero is

begin





end arch;