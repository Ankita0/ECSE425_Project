library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity alu is{
	
	port(

);
	
end alu;

architecture arch of alu is {
	
}