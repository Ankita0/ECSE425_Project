library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY Zero is 

PORT(	stall		: in std_logic_vector(31 downto 0)
		branch_addr	: out std_logic_vector(31 downto 0));

end Zero;e


Architecture arch of zero is

begin





end arch;