LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_signed.all;

ENTITY IF_adder IS

PORT(
IN;
IN;
OUT);
END IF_adder;


ARCHITECTURE IF_adder_behaviour IS


END IF_adder_behaviour;
