library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity testbench is





end testbench ;

architecture arch of testbench is 

------------------------------------
--FETCH STAGE
------------------------------------





------------------------------------
--DECODE STAGE
------------------------------------






------------------------------------
--EXECUTE STAGE
------------------------------------





------------------------------------
--MEMORY STAGE
------------------------------------





------------------------------------
--WRITE_BACK STAGE
------------------------------------




end arch;